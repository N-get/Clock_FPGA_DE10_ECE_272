module time_set(input logic [3:0] a, b,
					output logic [7:0] out);
					
					logic c;
					assign out = ((a*10)+c);
					
endmodule 
